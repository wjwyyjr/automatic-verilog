$header

// Local Variables:
// verilog-library-flags:("-f ../filelist/filelist.f")
// End:

`timescale 1ns/1ps

module $module_name
(
);
endmodule
